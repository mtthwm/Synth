module Synth (
	input wire clk,
	output wire gen_out
);

	assign gen_out = clk;

endmodule